module addr(parameter D=12)(
  
  
);