// Code your testbench here
// or browse Examples
`include "logical_sign_extend_tester.sv"