`include "logical_sign_extend.sv"